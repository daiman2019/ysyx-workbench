module data2seg(input[3:0] data,input neg_show,output [6:0] hout);
    reg [6:0] h;
    always @(*) begin
        case(data)//共阴极，输入为1对应数码管显示；若为共阳极，则对H取反
            4'b0000: h = 7'b0000000; // 0
            4'b0001: h = 7'b0000110; // 1
            4'b0010: h = 7'b1011011; // 2
            4'b0011: h = 7'b1001111; // 3
            4'b0100: h = 7'b0100110; // 4
            4'b0101: h = 7'b1101101; // 5
            4'b0110: h = 7'b1111101; // 6
            4'b0111: h = 7'b0000111; // 7
            4'b1000: h = 7'b1111111; // 8
            4'b1001: h = 7'b1101111; // 9
            4'b1010: h = 7'b1110111; // A
            4'b1011: h = 7'b1111100; // B
            4'b1100: h = 7'b0111001; // C
            4'b1101: h = 7'b1011110; // D
            4'b1110: h = 7'b1111001; // E
            4'b1111: h = 7'b1110001; // F
            default: h = 7'b0000000; // off
        endcase
    end
    assign hout = neg_show ? h : ~h; //共阴极，输入为1对应数码管显示；若为共阳极，则对H取反
endmodule


module key_identify(
    input clk,
    input resetn,
    input [7:0] data,
    output reg
)